----------------------------------------------------------------------------------------
-- Project       : RD53B Emulator
-- File          : rom_128x64bit_pkg.vhd
-- Description   : Expected output data from the model_yarr_rcv block in the RD53B testbench
-- Author        : gjones
----------------------------------------------------------------------------------------
library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

package rom_128x64bit_pkg is



--------------------------------------------------------------------------------
-- Expected output data from the model_yarr_rcv block in the RD53B testbench
--------------------------------------------------------------------------------
type     t_arr_hitdata_exp is array (0 to 127) of std_logic_vector(63 downto 0);
constant C_ARR_HITDATA_EXP   : t_arr_hitdata_exp := (
    X"8A10000100100002",    -- Tag = Tagbase 5 + 0
    X"0010000300100004",
    X"0010000500100006",
    X"0010000700100008",
    X"0020000100200002",
    X"0020000300200004",
    X"0020000500200006",
    X"0020000700200008",
    X"0030000100300002",
    X"0030000300300004",
    X"0030000500300006",
    X"0030000700300008",
    X"0040000100400002",
    X"0040000300400004",
    X"0040000500400006",
    X"0040000700400008",
    X"0050000100500002",
    X"0050000300500004",
    X"0050000500500006",
    X"005E0F07005E0F08",

    X"8A90000100100002",        -- Tagbase 5 + 1
    X"0010000300100004",
    X"0010000500100006",
    X"0010000700100008",
    X"0020000100200002",
    X"0020000300200004",
    X"0020000500200006",
    X"0020000700200008",
    X"0030000100300002",
    X"0030000300300004",
    X"0030000500300006",
    X"0030000700300008",
    X"0040000100400002",
    X"0040000300400004",
    X"0040000500400006",
    X"0040000700400008",
    X"0050000100500002",
    X"0050000300500004",
    X"0050000500500006",
    X"005E0F07005E0F08",

    X"8B10000100100002",        -- Tagbase 5 + 2
    X"0010000300100004",
    X"0010000500100006",
    X"0010000700100008",
    X"0020000100200002",
    X"0020000300200004",
    X"0020000500200006",
    X"0020000700200008",
    X"0030000100300002",
    X"0030000300300004",
    X"0030000500300006",
    X"0030000700300008",
    X"0040000100400002",
    X"0040000300400004",
    X"0040000500400006",
    X"0040000700400008",
    X"0050000100500002",
    X"0050000300500004",
    X"0050000500500006",
    X"005E0F07005E0F08",

    X"8B90000100100002",        -- Tagbase 5 + 3
    X"0010000300100004",
    X"0010000500100006",
    X"0010000700100008",
    X"0020000100200002",
    X"0020000300200004",
    X"0020000500200006",
    X"0020000700200008",
    X"0030000100300002",
    X"0030000300300004",
    X"0030000500300006",
    X"0030000700300008",
    X"0040000100400002",
    X"0040000300400004",
    X"0040000500400006",
    X"0040000700400008",
    X"0050000100500002",
    X"0050000300500004",
    X"0050000500500006",
    X"005E0F07005E0F08",

    X"8010000100100002",        -- Tagbase 0
    X"0010000300100004",
    X"0010000500100006",
    X"0010000700100008",
    X"0020000100200002",
    X"0020000300200004",
    X"0020000500200006",
    X"0020000700200008",
    X"0030000100300002",
    X"0030000300300004",
    X"0030000500300006",
    X"0030000700300008",
    X"0040000100400002",
    X"0040000300400004",
    X"0040000500400006",
    X"0040000700400008",
    X"0050000100500002",
    X"0050000300500004",
    X"0050000500500006",
    X"005E0F07005E0F08",

    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000",
    X"0000000000000000"
);
    
--type     t_arr_hitdata_exp is array (0 to 127) of std_logic_vector(63 downto 0);
--constant C_ARR_HITDATA_EXP   : t_arr_hitdata_exp := (
--    X"808300d5ff800000", 
--    X"0000000000000001", 
--    X"0000000000000002", 
--    X"0000000000000003", 
--    X"0000000000000004", 
--    X"0000000000000005", 
--    X"0000000000000006", 
--    X"0000000000000007", 
--    X"0000000000000008", 
--    X"0000000000000009", 
--    X"000000000000000A", 
--    X"000000000000000B", 
--    X"000000000000000C", 
--    X"000000000000000D", 
--    X"000000000000000E", 
--    X"000000000000000F", 
--    X"0000000000000010", 
--    X"0000000000000011", 
--    X"0000000000000012", 
--    X"0000000000000013", 
--    X"0000000000000014", 
--    X"0000000000000015", 
--    X"0000000000000016", 
--    X"0000000000000017", 
--    X"0000000000000018", 
--    X"0000000000000019", 
--    X"000000000000001A", 
--    X"000000000000001B", 
--    X"000000000000001C", 
--    X"000000000000001D", 
--    X"000000000000001E", 
--    X"000000000000001F", 
--    X"0000000000000020", 
--    X"0000000000000021", 
--    X"0000000000000022", 
--    X"0000000000000023", 
--    X"0000000000000024", 
--    X"0000000000000025", 
--    X"0000000000000026", 
--    X"0000000000000027", 
--    X"0000000000000028", 
--    X"0000000000000029", 
--    X"000000000000002A", 
--    X"000000000000002B", 
--    X"000000000000002C", 
--    X"000000000000002D", 
--    X"000000000000002E", 
--    X"000000000000002F", 
--    X"0000000000000030", 
--    X"0000000000000031", 
--    X"0000000000000032", 
--    X"0000000000000033", 
--    X"0000000000000034", 
--    X"0000000000000035", 
--    X"0000000000000036", 
--    X"0000000000000037", 
--    X"0000000000000038", 
--    X"0000000000000039", 
--    X"000000000000003A", 
--    X"000000000000003B", 
--    X"000000000000003C", 
--    X"000000000000003D", 
--    X"000000000000003E", 
--    X"000000000000003F", 
--    X"0000000000000040", 
--    X"0000000000000041", 
--    X"0000000000000042", 
--    X"0000000000000043", 
--    X"0000000000000044", 
--    X"0000000000000045", 
--    X"0000000000000046", 
--    X"0000000000000047", 
--    X"0000000000000048", 
--    X"0000000000000049", 
--    X"000000000000004A", 
--    X"000000000000004B", 
--    X"000000000000004C", 
--    X"000000000000004D", 
--    X"000000000000004E", 
--    X"000000000000004F", 
--    X"0000000000000050", 
--    X"0000000000000051", 
--    X"0000000000000052", 
--    X"0000000000000053", 
--    X"0000000000000054", 
--    X"0000000000000055", 
--    X"0000000000000056", 
--    X"0000000000000057", 
--    X"0000000000000058", 
--    X"0000000000000059", 
--    X"000000000000005A", 
--    X"000000000000005B", 
--    X"000000000000005C", 
--    X"000000000000005D", 
--    X"000000000000005E", 
--    X"000000000000005F", 
--    X"0000000000000060", 
--    X"0000000000000061", 
--    X"0000000000000062", 
--    X"0000000000000063", 
--    X"0000000000000064", 
--    X"0000000000000065", 
--    X"0000000000000066", 
--    X"0000000000000067", 
--    X"0000000000000068", 
--    X"0000000000000069", 
--    X"000000000000006A", 
--    X"000000000000006B", 
--    X"000000000000006C", 
--    X"000000000000006D", 
--    X"000000000000006E", 
--    X"000000000000006F", 
--    X"0000000000000070", 
--    X"0000000000000071", 
--    X"0000000000000072", 
--    X"0000000000000073", 
--    X"0000000000000074", 
--    X"0000000000000075", 
--    X"0000000000000076", 
--    X"0000000000000077", 
--    X"0000000000000078", 
--    X"0000000000000079", 
--    X"000000000000007A", 
--    X"000000000000007B", 
--    X"000000000000007C", 
--    X"000000000000007D", 
--    X"000000000000007E", 
--    X"000000000000007F" 
--);

end package rom_128x64bit_pkg;

















